// This module implements a working memory interface.
// It should be able to store message blocks in multiple locations.
// Ultimately it should indepenently load data while the hash function is running, reducing the
// amount of clock ticks necessary to generate a hash
module MOD_WORKING_MEM(CLK, D_IN, SLOT_ID, D_OUT );

output reg [31:0] OUT;
outpu 
input 
endmodule