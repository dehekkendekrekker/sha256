module MOD_EEPROM8K(
	input [0:12] A,
    output reg [0:7] IO,
	input CE,
	input OE,
	input WE
);

reg [0:7] buffer [0:8191];

initial begin
	// H constants
	buffer[0] = 8'h6a;
	buffer[1] = 8'h09;
	buffer[2] = 8'he6;
	buffer[3] = 8'h67;
	buffer[4] = 8'hbb;
	buffer[5] = 8'h67;
	buffer[6] = 8'hae;
	buffer[7] = 8'h85;
	buffer[8] = 8'h3c;
	buffer[9] = 8'h6e;
	buffer[10] = 8'hf3;
	buffer[11] = 8'h72;
	buffer[12] = 8'ha5;
	buffer[13] = 8'h4f;
	buffer[14] = 8'hf5;
	buffer[15] = 8'h3a;
	buffer[16] = 8'h51;
	buffer[17] = 8'h0e;
	buffer[18] = 8'h52;
	buffer[19] = 8'h7f;
	buffer[20] = 8'h9b;
	buffer[21] = 8'h05;
	buffer[22] = 8'h68;
	buffer[23] = 8'h8c;
	buffer[24] = 8'h1f;
	buffer[25] = 8'h83;
	buffer[26] = 8'hd9;
	buffer[27] = 8'hab;
	buffer[28] = 8'h5b;
	buffer[29] = 8'he0;
	buffer[30] = 8'hcd;
	buffer[31] = 8'h19;

	// K-Constants
	buffer[32] = 8'h42;
	buffer[33] = 8'h8a;
	buffer[34] = 8'h2f;
	buffer[35] = 8'h98;
	buffer[36] = 8'h71;
	buffer[37] = 8'h37;
	buffer[38] = 8'h44;
	buffer[39] = 8'h91;
	buffer[40] = 8'hb5;
	buffer[41] = 8'hc0;
	buffer[42] = 8'hfb;
	buffer[43] = 8'hcf;
	buffer[44] = 8'he9;
	buffer[45] = 8'hb5;
	buffer[46] = 8'hdb;
	buffer[47] = 8'ha5;
	buffer[48] = 8'h39;
	buffer[49] = 8'h56;
	buffer[50] = 8'hc2;
	buffer[51] = 8'h5b;
	buffer[52] = 8'h59;
	buffer[53] = 8'hf1;
	buffer[54] = 8'h11;
	buffer[55] = 8'hf1;
	buffer[56] = 8'h92;
	buffer[57] = 8'h3f;
	buffer[58] = 8'h82;
	buffer[59] = 8'ha4;
	buffer[60] = 8'hab;
	buffer[61] = 8'h1c;
	buffer[62] = 8'h5e;
	buffer[63] = 8'hd5;
	buffer[64] = 8'hd8;
	buffer[65] = 8'h07;
	buffer[66] = 8'haa;
	buffer[67] = 8'h98;
	buffer[68] = 8'h12;
	buffer[69] = 8'h83;
	buffer[70] = 8'h5b;
	buffer[71] = 8'h01;
	buffer[72] = 8'h24;
	buffer[73] = 8'h31;
	buffer[74] = 8'h85;
	buffer[75] = 8'hbe;
	buffer[76] = 8'h55;
	buffer[77] = 8'h0c;
	buffer[78] = 8'h7d;
	buffer[79] = 8'hc3;
	buffer[80] = 8'h72;
	buffer[81] = 8'hbe;
	buffer[82] = 8'h5d;
	buffer[83] = 8'h74;
	buffer[84] = 8'h80;
	buffer[85] = 8'hde;
	buffer[86] = 8'hb1;
	buffer[87] = 8'hfe;
	buffer[88] = 8'h9b;
	buffer[89] = 8'hdc;
	buffer[90] = 8'h06;
	buffer[91] = 8'ha7;
	buffer[92] = 8'hc1;
	buffer[93] = 8'h9b;
	buffer[94] = 8'hf1;
	buffer[95] = 8'h74;
	buffer[96] = 8'he4;
	buffer[97] = 8'h9b;
	buffer[98] = 8'h69;
	buffer[99] = 8'hc1;
	buffer[100] = 8'hef;
	buffer[101] = 8'hbe;
	buffer[102] = 8'h47;
	buffer[103] = 8'h86;
	buffer[104] = 8'h0f;
	buffer[105] = 8'hc1;
	buffer[106] = 8'h9d;
	buffer[107] = 8'hc6;
	buffer[108] = 8'h24;
	buffer[109] = 8'h0c;
	buffer[110] = 8'ha1;
	buffer[111] = 8'hcc;
	buffer[112] = 8'h2d;
	buffer[113] = 8'he9;
	buffer[114] = 8'h2c;
	buffer[115] = 8'h6f;
	buffer[116] = 8'h4a;
	buffer[117] = 8'h74;
	buffer[118] = 8'h84;
	buffer[119] = 8'haa;
	buffer[120] = 8'h5c;
	buffer[121] = 8'hb0;
	buffer[122] = 8'ha9;
	buffer[123] = 8'hdc;
	buffer[124] = 8'h76;
	buffer[125] = 8'hf9;
	buffer[126] = 8'h88;
	buffer[127] = 8'hda;
	buffer[128] = 8'h98;
	buffer[129] = 8'h3e;
	buffer[130] = 8'h51;
	buffer[131] = 8'h52;
	buffer[132] = 8'ha8;
	buffer[133] = 8'h31;
	buffer[134] = 8'hc6;
	buffer[135] = 8'h6d;
	buffer[136] = 8'hb0;
	buffer[137] = 8'h03;
	buffer[138] = 8'h27;
	buffer[139] = 8'hc8;
	buffer[140] = 8'hbf;
	buffer[141] = 8'h59;
	buffer[142] = 8'h7f;
	buffer[143] = 8'hc7;
	buffer[144] = 8'hc6;
	buffer[145] = 8'he0;
	buffer[146] = 8'h0b;
	buffer[147] = 8'hf3;
	buffer[148] = 8'hd5;
	buffer[149] = 8'ha7;
	buffer[150] = 8'h91;
	buffer[151] = 8'h47;
	buffer[152] = 8'h06;
	buffer[153] = 8'hca;
	buffer[154] = 8'h63;
	buffer[155] = 8'h51;
	buffer[156] = 8'h14;
	buffer[157] = 8'h29;
	buffer[158] = 8'h29;
	buffer[159] = 8'h67;
	buffer[160] = 8'h27;
	buffer[161] = 8'hb7;
	buffer[162] = 8'h0a;
	buffer[163] = 8'h85;
	buffer[164] = 8'h2e;
	buffer[165] = 8'h1b;
	buffer[166] = 8'h21;
	buffer[167] = 8'h38;
	buffer[168] = 8'h4d;
	buffer[169] = 8'h2c;
	buffer[170] = 8'h6d;
	buffer[171] = 8'hfc;
	buffer[172] = 8'h53;
	buffer[173] = 8'h38;
	buffer[174] = 8'h0d;
	buffer[175] = 8'h13;
	buffer[176] = 8'h65;
	buffer[177] = 8'h0a;
	buffer[178] = 8'h73;
	buffer[179] = 8'h54;
	buffer[180] = 8'h76;
	buffer[181] = 8'h6a;
	buffer[182] = 8'h0a;
	buffer[183] = 8'hbb;
	buffer[184] = 8'h81;
	buffer[185] = 8'hc2;
	buffer[186] = 8'hc9;
	buffer[187] = 8'h2e;
	buffer[188] = 8'h92;
	buffer[189] = 8'h72;
	buffer[190] = 8'h2c;
	buffer[191] = 8'h85;
	buffer[192] = 8'ha2;
	buffer[193] = 8'hbf;
	buffer[194] = 8'he8;
	buffer[195] = 8'ha1;
	buffer[196] = 8'ha8;
	buffer[197] = 8'h1a;
	buffer[198] = 8'h66;
	buffer[199] = 8'h4b;
	buffer[200] = 8'hc2;
	buffer[201] = 8'h4b;
	buffer[202] = 8'h8b;
	buffer[203] = 8'h70;
	buffer[204] = 8'hc7;
	buffer[205] = 8'h6c;
	buffer[206] = 8'h51;
	buffer[207] = 8'ha3;
	buffer[208] = 8'hd1;
	buffer[209] = 8'h92;
	buffer[210] = 8'he8;
	buffer[211] = 8'h19;
	buffer[212] = 8'hd6;
	buffer[213] = 8'h99;
	buffer[214] = 8'h06;
	buffer[215] = 8'h24;
	buffer[216] = 8'hf4;
	buffer[217] = 8'h0e;
	buffer[218] = 8'h35;
	buffer[219] = 8'h85;
	buffer[220] = 8'h10;
	buffer[221] = 8'h6a;
	buffer[222] = 8'ha0;
	buffer[223] = 8'h70;
	buffer[224] = 8'h19;
	buffer[225] = 8'ha4;
	buffer[226] = 8'hc1;
	buffer[227] = 8'h16;
	buffer[228] = 8'h1e;
	buffer[229] = 8'h37;
	buffer[230] = 8'h6c;
	buffer[231] = 8'h08;
	buffer[232] = 8'h27;
	buffer[233] = 8'h48;
	buffer[234] = 8'h77;
	buffer[235] = 8'h4c;
	buffer[236] = 8'h34;
	buffer[237] = 8'hb0;
	buffer[238] = 8'hbc;
	buffer[239] = 8'hb5;
	buffer[240] = 8'h39;
	buffer[241] = 8'h1c;
	buffer[242] = 8'h0c;
	buffer[243] = 8'hb3;
	buffer[244] = 8'h4e;
	buffer[245] = 8'hd8;
	buffer[246] = 8'haa;
	buffer[247] = 8'h4a;
	buffer[248] = 8'h5b;
	buffer[249] = 8'h9c;
	buffer[250] = 8'hca;
	buffer[251] = 8'h4f;
	buffer[252] = 8'h68;
	buffer[253] = 8'h2e;
	buffer[254] = 8'h6f;
	buffer[255] = 8'hf3;
	buffer[256] = 8'h74;
	buffer[257] = 8'h8f;
	buffer[258] = 8'h82;
	buffer[259] = 8'hee;
	buffer[260] = 8'h78;
	buffer[261] = 8'ha5;
	buffer[262] = 8'h63;
	buffer[263] = 8'h6f;
	buffer[264] = 8'h84;
	buffer[265] = 8'hc8;
	buffer[266] = 8'h78;
	buffer[267] = 8'h14;
	buffer[268] = 8'h8c;
	buffer[269] = 8'hc7;
	buffer[270] = 8'h02;
	buffer[271] = 8'h08;
	buffer[272] = 8'h90;
	buffer[273] = 8'hbe;
	buffer[274] = 8'hff;
	buffer[275] = 8'hfa;
	buffer[276] = 8'ha4;
	buffer[277] = 8'h50;
	buffer[278] = 8'h6c;
	buffer[279] = 8'heb;
	buffer[280] = 8'hbe;
	buffer[281] = 8'hf9;
	buffer[282] = 8'ha3;
	buffer[283] = 8'hf7;
	buffer[284] = 8'hc6;
	buffer[285] = 8'h71;
	buffer[286] = 8'h78;
	buffer[287] = 8'hf2;
end

always @* begin
	if (!CE && !OE && WE) begin
		IO <= buffer[A];
	end
end

endmodule

