module MOD_MAJORITY_TB;
`INIT

MOD_MAJORITY mut(
    E,F,G,Y
);

reg [0:31] E;
reg [0:31] F;
reg [0:31] G;
wire [0:31] Y;

localparam period = 20;  

initial begin
    `SET_MOD("MOD_MAJORITY_TB");
    $dumpfile("./build/MOD_MAJORITY_TB.vcd");
    $dumpvars(0, MOD_MAJORITY_TB);
    $timeformat(-6, 0, " us", 20);


    E = 32'b11111111111111111111111111111111; 
    F = 32'b11111111111111110000000000000000;
    G = 32'b11110000111100001111000011110000;
    #period
    if (Y != 32'b11111111111111111111000011110000)
        `FAILED("Test 1 failed");
    

    E = 32'b11111111111111110000000000000000; 
    F = 32'b11110000111100001111000011110000;
    G = 32'b11001100110011001100110011001100;
    #period
    if (Y != 32'b11111100111111001100000011000000) 
        `FAILED("Test 2 failed");

    E = 32'b11110000111100001111000011110000;
    F = 32'b11111100011000000000001110011111;
    G = 32'b10100101101001011010010110100101;
    #period
    if (Y != 32'b11110100111000001010000110110101) 
        `FAILED("Test 3 failed");

    E = 32'b11001100110011001100110011001100;
    F = 32'b10101010101010101010101010101010;
    G = 32'b11111111111111110000000000000000;
    #period
    if (Y != 32'b11101110111011101000100010001000) 
        `FAILED("Test 4 failed");

    E = 32'b10101010101010101010101010101010;
    F = 32'b10100101101001011010010110100101;
    G = 32'b11111100011000000000001110011111;
    #period
    if (Y != 32'b10101100101000001010001110101111) 
        `FAILED("Test 5 failed");



  


end

endmodule