// This module ties everything together

`include "./src/verilog/MOD_COMPRESSOR.v"
module MOD_SHA256(CLK);

input CLK;

MOD_COMPRESSOR compressor(CLK, RESET, I, W, K, 
H[0],H[1],H[2],H[3],H[4],H[5],H[6],H[7],
R[0],R[1],R[2],R[3],R[4],R[5],R[6],R[7]);

// We should be some logic that copies the H values into the latches
// Latches should be implemented here

reg [31:0] H [8];
reg [31:0] R [8];

reg RESET;
reg [5:0] I;
reg [31:0] W, K;










endmodule



// // Letter registers
// reg [31:0] a;
// reg [31:0] b;
// reg [31:0] c;
// reg [31:0] d;
// reg [31:0] e;
// reg [31:0] f;
// reg [31:0] g;
// reg [31:0] h;
// reg [31:0] Temp1;
// reg [31:0] Temp2;


// reg [31:0] H [8];
// reg [31:0] W [128];





// initial begin
//     state = ST_IDLE;
//     ctr_clr = 1;


//     H[0] = 32'h6a09e667;
//     H[1] = 32'hbb67ae85;
//     H[2] = 32'h3c6ef372;
//     H[3] = 32'h54ff53a;
//     H[4] = 32'h10e527f;
//     H[5] = 32'h9b05688c;
//     H[6] = 32'h1f83d9ab;
//     H[7] = 32'h5be0cd19;

//     W[0] = 32'b01001000011001010110110001101100;
//     W[1] = 32'b01101111001000000111011101101111;
//     W[2] = 32'b01110010011011000110010000100001;
//     W[3] = 32'b10000000000000000000000000000000;
//     W[4] = 32'b00000000000000000000000000000000;
//     W[5] = 32'b00000000000000000000000000000000;
//     W[6] = 32'b00000000000000000000000000000000;
//     W[7] = 32'b00000000000000000000000000000000;
//     W[8] = 32'b00000000000000000000000000000000;
//     W[9] = 32'b00000000000000000000000000000000;
//     W[10] = 32'b00000000000000000000000000000000;
//     W[11] = 32'b00000000000000000000000000000000;
//     W[12] = 32'b00000000000000000000000000000000;
//     W[13] = 32'b00000000000000000000000000000000;
//     W[14] = 32'b00000000000000000000000000000000;
//     W[15] = 32'b00000000000000000000000001100000;

//     // TODO: Fill this with representative data
//     W[16] = 32'b00000000000000000000000000000000;
//     W[17] = 32'b00000000000000000000000000000000;
//     W[18] = 32'b00000000000000000000000000000000;
//     W[19] = 32'b00000000000000000000000000000000;
//     W[20] = 32'b00000000000000000000000000000000;
//     W[21] = 32'b00000000000000000000000000000000;
//     W[22] = 32'b00000000000000000000000000000000;
//     W[23] = 32'b00000000000000000000000000000000;
//     W[24] = 32'b00000000000000000000000000000000;
//     W[25] = 32'b00000000000000000000000000000000;
//     W[26] = 32'b00000000000000000000000000000000;
//     W[27] = 32'b00000000000000000000000000000000;
//     W[28] = 32'b00000000000000000000000000000000;
//     W[29] = 32'b00000000000000000000000000000000;
//     W[30] = 32'b00000000000000000000000000000000;
//     W[31] = 32'b00000000000000000000000000000000;

// end





// endmodule