`include "./src/verilog/7400/MOD_74x393.v"
`include "./src/verilog/MOD_S0.v"
`include "./src/verilog/MOD_S1.v"
module MOD_SHA256(
    input CLK,
    output [31:0] W_OUT
);

MOD_74x393 h_init_ctr(CLK,ctr_clr, hi[3],ctr_clr, hi[3:0], hi[7:4]);
MOD_S0 s0(s0_in, s0_out);
MOD_S1 s1(s1_in, s1_out);


reg [7:0] hi;
reg ctr_clr;

assign W_OUT = W[hi];

reg [31:0] s0_in, s0_out;
reg [31:0] s1_in, s1_out;


// Letter registers
reg [31:0] a;
reg [31:0] b;
reg [31:0] c;
reg [31:0] d;
reg [31:0] e;
reg [31:0] f;
reg [31:0] g;
reg [31:0] h;
reg [31:0] Temp1;
reg [31:0] Temp2;


reg [31:0] H [8];
reg [31:0] W [64];


reg [1:0] state;

localparam ST_IDLE = 0;
localparam ST_INIT = 1;
localparam ST_PROC_W = 2;
localparam ST_DONE = 3;

initial begin
    state = ST_IDLE;
    ctr_clr = 1;


    H[0] = 32'h6a09e667;
    H[1] = 32'hbb67ae85;
    H[2] = 32'h3c6ef372;
    H[3] = 32'h54ff53a;
    H[4] = 32'h10e527f;
    H[5] = 32'h9b05688c;
    H[6] = 32'h1f83d9ab;
    H[7] = 32'h5be0cd19;

    W[0] = 32'b01001000011001010110110001101100;
    W[1] = 32'b01101111001000000111011101101111;
    W[2] = 32'b01110010011011000110010000100001;
    W[3] = 32'b10000000000000000000000000000000;
    W[4] = 32'b00000000000000000000000000000000;
    W[5] = 32'b00000000000000000000000000000000;
    W[6] = 32'b00000000000000000000000000000000;
    W[7] = 32'b00000000000000000000000000000000;
    W[8] = 32'b00000000000000000000000000000000;
    W[9] = 32'b00000000000000000000000000000000;
    W[10] = 32'b00000000000000000000000000000000;
    W[11] = 32'b00000000000000000000000000000000;
    W[12] = 32'b00000000000000000000000000000000;
    W[13] = 32'b00000000000000000000000000000000;
    W[14] = 32'b00000000000000000000000000000000;
    W[15] = 32'b00000000000000000000000001100000;


    W[16] = 32'b00000000000000000000000000000000;
    W[17] = 32'b00000000000000000000000000000000;
    W[18] = 32'b00000000000000000000000000000000;
    W[19] = 32'b00000000000000000000000000000000;
    W[20] = 32'b00000000000000000000000000000000;
    W[21] = 32'b00000000000000000000000000000000;
    W[22] = 32'b00000000000000000000000000000000;
    W[23] = 32'b00000000000000000000000000000000;
    W[24] = 32'b00000000000000000000000000000000;
    W[25] = 32'b00000000000000000000000000000000;
    W[26] = 32'b00000000000000000000000000000000;
    W[27] = 32'b00000000000000000000000000000000;
    W[28] = 32'b00000000000000000000000000000000;
    W[29] = 32'b00000000000000000000000000000000;
    W[30] = 32'b00000000000000000000000000000000;
    W[31] = 32'b00000000000000000000000000000000;

    W[32] = 32'b00000000000000000000000000000000;
    W[33] = 32'b00000000000000000000000000000000;
    W[34] = 32'b00000000000000000000000000000000;
    W[35] = 32'b00000000000000000000000000000000;
    W[36] = 32'b00000000000000000000000000000000;
    W[37] = 32'b00000000000000000000000000000000;
    W[38] = 32'b00000000000000000000000000000000;
    W[39] = 32'b00000000000000000000000000000000;
    W[40] = 32'b00000000000000000000000000000000;
    W[41] = 32'b00000000000000000000000000000000;
    W[42] = 32'b00000000000000000000000000000000;
    W[43] = 32'b00000000000000000000000000000000;
    W[44] = 32'b00000000000000000000000000000000;
    W[45] = 32'b00000000000000000000000000000000;
    W[46] = 32'b00000000000000000000000000000000;
    W[47] = 32'b00000000000000000000000000000000;

    W[48] = 32'b00000000000000000000000000000000;
    W[49] = 32'b00000000000000000000000000000000;
    W[50] = 32'b00000000000000000000000000000000;
    W[51] = 32'b00000000000000000000000000000000;
    W[52] = 32'b00000000000000000000000000000000;
    W[53] = 32'b00000000000000000000000000000000;
    W[54] = 32'b00000000000000000000000000000000;
    W[55] = 32'b00000000000000000000000000000000;
    W[56] = 32'b00000000000000000000000000000000;
    W[57] = 32'b00000000000000000000000000000000;
    W[58] = 32'b00000000000000000000000000000000;
    W[59] = 32'b00000000000000000000000000000000;
    W[60] = 32'b00000000000000000000000000000000;
    W[61] = 32'b00000000000000000000000000000000;
    W[62] = 32'b00000000000000000000000000000000;
    W[63] = 32'b00000000000000000000000000000000;
end



always @(negedge CLK) begin
    if (state == ST_IDLE) begin
        state <= ST_INIT;
    end
    


end

always @(posedge CLK) begin
    if (state == ST_PROC_W) begin
        s0_in <= W[hi + 1];
        s1_in <= W[hi + 14];
    end
end


reg [31:0] w0, w9;

assign w0 = W[hi];

always @(negedge CLK) begin
    if (state == ST_PROC_W) begin
        $display("i: %d s0_in: %b s0_out: %b", hi, s0_in,s0_out);
        //$display("s1_out: %b", s1_out);


        w0 = W[hi];
        w9 = W[hi + 9];
        


        W[hi + 16] <= w0 + s0_out + w9 + s1_out;

        

        if (hi == 48) begin
            state <= ST_DONE;
        end

    end
end



always @(state) begin
    if (state == ST_INIT) begin
        a <= H[0];
        b <= H[1];
        c <= H[2];
        d <= H[3];
        e <= H[4];
        f <= H[5];
        g <= H[6];
        h <= H[7];
        Temp1 <= 0;
        Temp2 <= 1;

        ctr_clr <= 0;
        state <= ST_PROC_W;
    end
end


endmodule