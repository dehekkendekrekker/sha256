module MOD_CHOICE_TB;
`INIT

MOD_CHOICE mut(
    E,F,G,Y
);

reg [0:31] E;
reg [0:31] F;
reg [0:31] G;
wire [0:31] Y;

localparam period = 20;  

initial begin
    `SET_MOD("MOD_CHOICE_TB");
    $dumpfile("./build/MOD_CHOICE_TB.vcd");
    $dumpvars(0, MOD_CHOICE_TB);
    $timeformat(-6, 0, " us", 20);


    E = 32'b11111111111111111111111111111111; 
    F = 32'b11111111111111110000000000000000;
    G = 32'b11110000111100001111000011110000;
    #period
    if (Y != 32'b11111111111111110000000000000000)
        `FAILED("Test 1 failed");
    

    E = 32'b11111111111111110000000000000000; 
    F = 32'b11110000111100001111000011110000;
    G = 32'b11001100110011001100110011001100;
    #period
    if (Y != 32'b11110000111100001100110011001100) 
        `FAILED("Test 2 failed");

    E = 32'b11110000111100001111000011110000;
    F = 32'b11111100011000000000001110011111;
    G = 32'b10100101101001011010010110100101;
    #period
    if (Y != 32'b11110101011001010000010110010101) 
        `FAILED("Test 3 failed");

    E = 32'b11001100110011001100110011001100;
    F = 32'b10101010101010101010101010101010;
    G = 32'b11111111111111110000000000000000;
    #period
    if (Y != 32'b10111011101110111000100010001000) 
        `FAILED("Test 4 failed");

    E = 32'b10101010101010101010101010101010;
    F = 32'b10100101101001011010010110100101;
    G = 32'b11111100011000000000001110011111;
    #period
    if (Y != 32'b11110100111000001010000110110101) 
        `FAILED("Test 5 failed");



  


end

endmodule