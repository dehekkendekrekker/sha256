module MOD_EEPROM8K_1 (A, IO, CE, OE, WE); 

input [0:12] A;
inout [0:7] IO;
input CE;
input OE;
input WE;

MOD_EEPROM8K __TECHMAP_REPLACE_ (.A(A), .IO(IO), .CE(CE), .OE(OE), .WE(WE)); 

endmodule

module MOD_EEPROM8K_2 (A, IO, CE, OE, WE); 

input [0:12] A;
inout [0:7] IO;
input CE;
input OE;
input WE;

MOD_EEPROM8K __TECHMAP_REPLACE_ (.A(A), .IO(IO), .CE(CE), .OE(OE), .WE(WE)); 

endmodule

module MOD_EEPROM8K_3 (A, IO, CE, OE, WE); 

input [0:12] A;
inout [0:7] IO;
input CE;
input OE;
input WE;

MOD_EEPROM8K __TECHMAP_REPLACE_ (.A(A), .IO(IO), .CE(CE), .OE(OE), .WE(WE)); 

endmodule

module MOD_EEPROM8K_4 (A, IO, CE, OE, WE); 

input [0:12] A;
inout [0:7] IO;
input CE;
input OE;
input WE;

MOD_EEPROM8K __TECHMAP_REPLACE_ (.A(A), .IO(IO), .CE(CE), .OE(OE), .WE(WE)); 

endmodule